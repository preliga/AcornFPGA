----------------------------------
-- Łukasz DZIEŁ (883533374)     --
-- FPGACOMMEXAMPLE-v2           --
-- 01.2016                      --
-- 1.0                          --
----------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY memory IS PORT
(	
	CLK		:IN STD_LOGIC;
	
	DIN	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	ADDR_RD	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	RD   		:IN STD_LOGIC;
	
	ADDR_WR	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	WR			:IN STD_LOGIC;
	
	DOUT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE A1 OF memory IS
	TYPE MEMORY_BLOCK IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEM : MEMORY_BLOCK;
BEGIN
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (WR = '1') THEN
				MEM(conv_integer(ADDR_WR)) <= DIN;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF(RD = '1') THEN
				DOUT <= MEM(conv_integer(ADDR_RD));
			ELSE
				DOUT <= (others => '0');
			END IF;
		END IF;
	END PROCESS;
	
END ARCHITECTURE;