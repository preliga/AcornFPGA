LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY m IS PORT
(
	INP	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	KEY_S	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	OPT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE A1 OF m IS
BEGIN
	OPT <= INP xor KEY_S;
END ARCHITECTURE;