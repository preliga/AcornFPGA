LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY status_multiplexer IS PORT
(
	DATA_INP		:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	--STATUS		:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	WR_STATUS	:IN STD_LOGIC_vector(1 downto 0);
	
	DATA_OPT		:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE A1 OF status_multiplexer IS
BEGIN
	WITH WR_STATUS SELECT
		DATA_OPT <= DATA_INP 						WHEN "11",
					(30 downto 0 =>'0', 31 =>'1')	WHEN "01",
					(31 downto 0 =>'0')				WHEN others;
END ARCHITECTURE;