LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FBK128 IS PORT
(
	S		:IN STD_LOGIC_VECTOR(292 downto 0);
	KS		:IN STD_LOGIC_VECTOR(31 downto 0);
	CA		:IN STD_LOGIC;
	CB		:IN STD_LOGIC;
	
	OPT	:OUT STD_LOGIC_VECTOR(31 downto 0)
);
END ENTITY;

ARCHITECTURE A1 OF FBK128 IS
BEGIN
END ARCHITECTURE;