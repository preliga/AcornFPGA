LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY key IS PORT
(
	CLK	:IN STD_LOGIC;
	
	RD		:IN STD_LOGIC;
	WR		:IN STD_LOGIC;
	
	ADR	:IN STD_LOGIC_VECTOR(1 downto 0);
	INP	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	OPT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE A1 OF key IS
	TYPE MEM_REGISTER IS ARRAY (0 TO 3) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL KEY_REGISTER : MEM_REGISTER;
BEGIN

	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (WR = '1') THEN
				KEY_REGISTER(conv_integer(ADR)) <= INP;
			END IF;
		END IF;
	END PROCESS;

	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (RD = '1') THEN
				OPT <= KEY_REGISTER(conv_integer(ADR));
			END IF;
		END IF;
	END PROCESS;
	
END ARCHITECTURE;