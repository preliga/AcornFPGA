LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY state IS PORT
(
	CLK	:IN STD_LOGIC;
	INP_F	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	INP_M	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	WR		:IN STD_LOGIC;
	RESET	:IN STD_LOGIC;
	S		:OUT STD_LOGIC_VECTOR(292 downto 0)
);
END ENTITY;

ARCHITECTURE A1 OF state IS
	SIGNAL STATE : STD_LOGIC_VECTOR(292 DOWNTO 0);
	
BEGIN

	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (WR = '1') THEN
				
				STATE <= (INP_M XOR INP_F) & STATE(292 downto 32);
				
				
				
			END IF;
		END IF;
	END PROCESS;
	
	S <= STATE;
	
END ARCHITECTURE;