LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY add_one IS PORT
(
	DATA_INP	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	ADD_ONE	:IN STD_LOGIC;
	
	DATA_OPT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE A1 OF add_one IS
BEGIN
	DATA_OPT <= (DATA_INP(0) xor ADD_ONE) & DATA_INP(31 downto 1);
END ARCHITECTURE;