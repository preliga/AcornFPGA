----------------------------------
-- Łukasz DZIEŁ (883533374)     --
-- FPGACOMMEXAMPLE-v2           --
-- 01.2016                      --
-- 1.0                          --
----------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY WORK;
USE WORK.ALL;
USE WORK.RS232_INTERFACE_PKG.ALL;

ENTITY RS232_TRANSMITTER IS PORT
(	
	CLK	:IN STD_LOGIC;
	INIT	:IN STD_LOGIC;
	DRL	:IN STD_LOGIC;
	LOAD	:OUT STD_LOGIC;
	DIN	:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	TX		:OUT STD_LOGIC
);
END ENTITY;

ARCHITECTURE RS232_RS232_TRANSMITTER OF RS232_TRANSMITTER IS
	
	SIGNAL FSM 						:STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL BIT_COUNTER 			:STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL CLOCK_COUNTER 		:STD_LOGIC_VECTOR(15 DOWNTO 0); 	
	SIGNAL TRANSMIT_REGISTER 	:STD_LOGIC_VECTOR(9 DOWNTO 0);
	SIGNAL TX_REG 					:STD_LOGIC := '1';
	
BEGIN

	PROCESS(CLK, INIT)
	BEGIN
		IF (INIT = '1') THEN FSM <= X"0";
		ELSIF(CLK'EVENT AND CLK = '1') THEN
			CASE FSM IS
				WHEN X"0" =>	IF(DRL = '1') THEN
										FSM <= X"1";
									END IF;
				
				WHEN X"1" =>	FSM <= X"2";
				WHEN X"2" =>	FSM <= X"3";
				WHEN X"3" =>	FSM <= X"4";
				WHEN X"4" =>	IF(CLOCK_COUNTER = X"0000") THEN
										FSM <= X"5"; 
									END IF;	
				WHEN X"5" => 	IF(BIT_COUNTER = X"0")THEN
										FSM <= X"0";
									ELSE
										FSM <= X"3";
									END IF;
				WHEN OTHERS => FSM <= X"0";						
			END CASE;
		END IF;
	END PROCESS;


	PROCESS(CLK, INIT)
	BEGIN
		IF(INIT = '1') THEN BIT_COUNTER <= (others => '0');
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			IF(FSM = X"2") THEN
				BIT_COUNTER <= X"A";
			END IF;
			IF(FSM = X"3") THEN
				BIT_COUNTER <= STD_LOGIC_VECTOR(unsigned(BIT_COUNTER) - 1);
			END IF;
		END IF;
	END PROCESS;

	PROCESS(CLK, INIT)
	BEGIN
		IF(INIT = '1') THEN CLOCK_COUNTER <= (others => '0');
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			IF(FSM = X"3") THEN
				CLOCK_COUNTER <= BIT_RATE_VAL;
			END IF;
			IF(FSM = X"4") THEN
				CLOCK_COUNTER <= STD_LOGIC_VECTOR(unsigned(CLOCK_COUNTER) - 1);
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CLK, INIT)
	BEGIN
		IF(INIT = '1') THEN TRANSMIT_REGISTER <= "0000000000";
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			IF(FSM = X"2") THEN
				TRANSMIT_REGISTER <= '1' & DIN & '0';
			END IF;
			IF(FSM = X"3") THEN
				TRANSMIT_REGISTER <= '0' & TRANSMIT_REGISTER(9 DOWNTO 1);
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CLK, INIT)
	BEGIN
		IF(INIT = '1') THEN TX_REG <= '1';
		ELSIF(CLK'EVENT AND CLK = '1') THEN
			IF(FSM = X"3") THEN
				TX_REG <= TRANSMIT_REGISTER(0);
			END IF;
		END IF;
	END PROCESS;
	
	LOAD	<= '1' WHEN FSM = X"1" ELSE '0';
	TX		<= TX_REG;
	
END ARCHITECTURE;