LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY token_checker IS PORT
(
	DATA_IN	:IN STD_LOGIC_VECTOR(31 downto 0);
	IS_ZERO	:OUT STD_LOGIC
);
END ENTITY;

ARCHITECTURE A1 OF token_checker IS
BEGIN
	IS_ZERO <= 	DATA_IN(0) OR DATA_IN(1) OR DATA_IN(2) OR DATA_IN(3) OR
					DATA_IN(4) OR DATA_IN(5) OR DATA_IN(6) OR DATA_IN(7) OR
					DATA_IN(8) OR DATA_IN(9) OR DATA_IN(10) OR DATA_IN(11) OR
					DATA_IN(12) OR DATA_IN(13) OR DATA_IN(14) OR DATA_IN(15) OR
					DATA_IN(16) OR DATA_IN(17) OR DATA_IN(18) OR DATA_IN(19) OR
					DATA_IN(20) OR DATA_IN(21) OR DATA_IN(22) OR DATA_IN(23) OR
					DATA_IN(24) OR DATA_IN(25) OR DATA_IN(26) OR DATA_IN(27) OR
					DATA_IN(28) OR DATA_IN(29) OR	DATA_IN(30) OR DATA_IN(31);
END ARCHITECTURE;